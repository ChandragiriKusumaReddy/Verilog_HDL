module mux_16x1(
  input [15:0] i,
  input [3:0] s,
  output y );
  assign y = (~s[3]&~s[2]&~s[1]&~s[0]&i[0]) |
    (~s[3]&~s[2]&~s[1]&s[0]&i[1]) |
    (~s[3]&~s[2]&s[1]&~s[0]&i[2]) |
    (~s[3]&~s[2]&s[1]&s[0]&i[3])  |
    (~s[3]&s[2]&~s[1]&~s[0]&i[4]) |
    (~s[3]&s[2]&~s[1]&s[0]&i[5])  |
    (~s[3]&s[2]&s[1]&~s[0]&i[6])  |
    (~s[3]&s[2]&s[1]&s[0]&i[7])   |
    (s[3]&~s[2]&~s[1]&~s[0]&i[8]) |
    (s[3]&~s[2]&~s[1]&s[0]&i[9])  |
    (s[3]&~s[2]&s[1]&~s[0]&i[10]) |
    (s[3]&~s[2]&s[1]&s[0]&i[11])  |
    (s[3]&s[2]&~s[1]&s~[0]&i[12]) |
    (s[3]&s[2]&~s[1]&s[0]&i[13])  |
    (s[3]&s[2]&s[1]&~s[0]&i[14])  |
    (s[3]&s[2]&s[1]&s[0]&i[15]) ;
endmodule
